* Extracted by KLayout with SG13G2 LVS runset on : 28/04/2025 03:36

.SUBCKT TOP \$3.VBB2 \$3.VBB1
C$1 \$I3 \$1 cap_cmim w=20u l=25u A=500p P=90u m=8
C$4 \$3.VBB1 \$1 cap_cmim w=20u l=25u A=500p P=90u m=6
C$10 \$3.VBB2 \$1 cap_cmim w=20u l=25u A=500p P=90u m=4
R$19 \$I27 \$3.VBB2 rhigh w=2u l=5.5u ps=0 b=0 m=1
R$20 \$I28 \$I3 rsil w=7.5u l=5.5u ps=0 b=0 m=1
Q$21 \$I28 \$I27 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=12.988p PB=15.62u
+ AC=12.976684p PC=15.61u NE=2 m=2
Q$23 \$I25 \$I26 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=12.988p PB=15.62u
+ AC=12.976684p PC=15.61u NE=2 m=2
R$25 \$I26 \$3.VBB1 rhigh w=1.9u l=5.5u ps=0 b=0 m=1
R$26 \$I23 \$3.VBB1 rhigh w=1.9u l=5.5u ps=0 b=0 m=1
R$27 \$I25 \$I3 rsil w=7.5u l=5u ps=0 b=0 m=1
R$28 \$I24 \$I3 rsil w=7.5u l=5u ps=0 b=0 m=1
R$29 \$I21 \$I3 rsil w=7.5u l=5u ps=0 b=0 m=1
Q$30 \$I24 \$I23 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=25.605p PB=23.02u
+ AC=25.589984p PC=23.01u NE=4 m=4
Q$34 \$I21 \$I22 \$1 \$1 npn13G2 AE=0.063p PE=1.94u AB=25.605p PB=23.02u
+ AC=25.589984p PC=23.01u NE=4 m=4
R$38 \$I22 \$3.VBB1 rhigh w=1.9u l=7u ps=0 b=0 m=1
.ENDS TOP
